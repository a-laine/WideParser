


/*
	Class Description Language :
	
	+ les accolades {} définissent une classe d'association (map)
	  où chaques paire est notée:  clée : valeur
	+ les crochets [] définissent un conteneur à valeur indicée
	+ les , ou ; délimitent les éléments dans les types composés
	+ types primitifs (ou scalaires):
		- booléen
		- entier
		- réel
		- chaine de caractères, sont délimitées par '' ou "", "" gère les échappements
		  une chaine de 1 caractère est considéré comme un caractère plutot
		  que comme une chaine
	+ toute variable peut être renseignée par un nom lorsqu'elle est déclaré dans la racine
	  elle est alors suivie par un signe = ou :
	+ un nom de variable ou la clé d'une classe d'association peut contenir des caractères
	  spéciaux en l'écrivant comme une chaine de caractère, donc avec '' ou "", sinon elle doit être
	  uniquement composés de caractères alphanumériques et comencer par une lettre
	  la notation "" permet l'echappement de caractères
	+ une variable nomée peut être référencé plus tard dans le code en suffixant son nom par @
*/




//Définition d' une classe d'association globale
myClass :
{
	id : "myObject",	#une chaine
	att1 : true,		#constante
	att2 : 150,			#nombre
	att3 : @unObjet,	#une référence
	att4 : [10, 25, 6],	#un tableau
	att5 : {1:'a', 2:'b', 3:'c'}, #une "map"
}